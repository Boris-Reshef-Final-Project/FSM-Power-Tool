library ieee;
use ieee.std_logic_1164.all;

package tb_package_$ is

  -- constants and types
  constant num_inputs   : positive  := ?x; -- number of inputs
  constant num_outputs  : positive  := ?y; -- number of outputs
  constant num_clocks   : positive  := ?c; -- number of clocks
  constant clk_period   : time      := ?p;
  -- state type
  ?s
    
  -- file names and locations
  constant kis_src_path : string    := ?k; -- file path of source .kis file

end package tb_package_$;


package body tb_package_$ is
end package body tb_package_$;