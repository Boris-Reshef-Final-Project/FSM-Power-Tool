library ieee;
use ieee.std_logic_1164.all;

package $_tb_pack is

  -- constants and types
  constant num_inputs   : positive  := ~;
  constant num_outputs  : positive  := ~;
  constant num_clocks   : positive  := ~;
  constant clk_freq     : positive  := ~; -- in MHz  
  constant clk_period   : time      := ~ ns;
  type state is (~);
    
  -- file names and locations
  constant kis_src_path : string    := ~; -- file path of source .kis file

end package $_tb_pack;


package body $_tb_pack is
end package body $_tb_pack;