Library IEEE;
use ieee.std_logic_1164.all;
library work;
use work.all;
use work.top_pack_$.all;
library altera; 
use altera.altera_primitives_components.all;
library altera_mf;
use altera_mf.altera_mf_components.all;
library cycloneive_atoms;
use cycloneive_atoms.all;
library cycloneive_components;
use cycloneive_components.all;

entity top_$ is
    generic (
        simulation_mode : boolean := false;
        power_analyzer  : boolean := true;
        baseline_power  : boolean := false;
        full_fpga       : boolean := false;
        duplicates      : integer := 100
    );
    port(
        rst	    : in	std_logic := '1';
        clk	: in    std_logic;
        x		: in	std_logic_vector(?x downto 0) := (others => '0');
        y		: out	std_logic_vector(?y downto 0) := (others => '0')	
    );
    -- Connect the pins to the FPGA for tests on the board
    attribute altera_chip_pin_lc              : string;
    attribute altera_chip_pin_lc of clk       : signal is "Y2";     -- 50 MHz clock from the board
    attribute altera_chip_pin_lc of rst       : signal is "AB28";   -- Reset switch: Slide switch 0

    end entity top_$;
 
    
architecture arc_top of top_$ is
    
        signal clken, clk_out, S, PLL_clk	: std_logic_vector(?c downto 0) := (0 => '1', others => '0');
        signal LFSR_out  : std_logic_vector(x'range) := (others => '1');
        signal fsm_input : std_logic_vector(x'range) := (others => '0');
    
    begin

        -- when working in software, the inputs are generated by the software
        -- but when working in the hardware (on the board), the inputs are generated by an LFSR
        fsm_input <= LFSR_out when (baseline_power or full_fpga) else x;

        -- generate 1 FSM
        -- Used in: simulation, power analyzer, full_fpga
        G_FSM: if (not baseline_power) generate
            FSM: entity work.$
            port map(
                rst	    => rst,
                clk	    => clk_out,
                x		=> fsm_input,
                y		=> y,
                clken	=> clken
                );
        end generate G_FSM;


        -- generate many FSMs to fill the area on the chip to about 30%
        -- change the value of 'duplicates' (generic) to control the amount of FSMs
        -- Used in: power_analyzer, full_fpga
        G_MANY_FSMS: if (full_fpga or power_analyzer) generate
            G_FSM_LOOP: for i in 0 to duplicates generate
                FSM_area_fill: entity work.$
                    port map(
                        rst	    => rst,
                        clk	    => clk_out,
                        x		=> fsm_input,
                        y		=> open,
                        clken	=> open
                        );
            end generate G_FSM_LOOP;
            
        end generate G_MANY_FSMS;

        -- generate PLLs
        -- Used in: simulation, power_analyzer, full_fpga
        G_PLL: if not baseline_power generate
            G_PLL_LOOP: for i in 0 to ?c generate
                PLL: PLL_altpll PORT MAP (
                    inclk0  => clk,
                    clken   => clken(i),
                    clk_out => clk_out(i)
                );
            end generate G_PLL_LOOP;
        end generate G_PLL;

        -- generate LFSR
        -- Used in: baseline_power, full_fpga
        G_LFSR: if (baseline_power or full_fpga) generate
            process(clk) is
            begin
                if (rst = '1') then
                    LFSR_out <= (others => '1');
                elsif rising_edge(clk) then
                    LFSR_out <= LFSR(LFSR_out, c_polynom);
                    if (baseline_power) then -- to make sure the LFSR is actually driving something
                        fsm_input <= y;
                    end if;
                end if;
            end process;
        end generate G_LFSR;
         
end architecture arc_top;